$date
	Tue Jul 28 20:53:00 2020
$end
$version
	Icarus Verilog
$end
$timescale
	1ns
$end
$scope module osl_tb $end
$var wire 32 ! hostB_dout_w [31:0] $end
$var wire 1 " hostB_dor_w $end
$var wire 1 # hostB_dir_w $end
$var wire 32 $ hostA_dout_w [31:0] $end
$var wire 1 % hostA_dor_w $end
$var wire 1 & hostA_dir_w $end
$var wire 1 ' data1_w $end
$var wire 1 ( data0_w $end
$var reg 1 ) clk_r $end
$var reg 32 * hostA_din_r [31:0] $end
$var reg 1 + hostA_rd_r $end
$var reg 1 , hostA_wr_r $end
$var reg 32 - hostB_din_r [31:0] $end
$var reg 1 . hostB_rd_r $end
$var reg 1 / hostB_wr_r $end
$var reg 1 0 rstb_r $end
$var reg 1 1 tx_r $end
$scope module UA_0 $end
$var wire 1 ) clk $end
$var wire 2 2 din_w [1:0] $end
$var wire 32 3 host_din [31:0] $end
$var wire 32 4 host_dout [31:0] $end
$var wire 1 + host_rd $end
$var wire 1 , host_wr $end
$var wire 1 0 resetb $end
$var wire 1 ' tx $end
$var wire 1 ( rx $end
$var wire 1 % host_dor $end
$var wire 1 & host_dir $end
$var reg 2 5 din_q [1:0] $end
$var reg 32 6 par2ser_q [31:0] $end
$var reg 1 7 rx_ack_req_q $end
$var reg 5 8 rx_count_q [4:0] $end
$var reg 1 9 rx_ready_q $end
$var reg 2 : rx_state_q [1:0] $end
$var reg 32 ; ser2par_q [31:0] $end
$var reg 1 < tx_ack_rcvd_q $end
$var reg 5 = tx_count_q [4:0] $end
$var reg 1 > tx_r $end
$var reg 1 ? tx_ready_q $end
$var reg 3 @ tx_state_q [2:0] $end
$upscope $end
$scope module UB_1 $end
$var wire 1 ) clk $end
$var wire 2 A din_w [1:0] $end
$var wire 32 B host_din [31:0] $end
$var wire 32 C host_dout [31:0] $end
$var wire 1 . host_rd $end
$var wire 1 / host_wr $end
$var wire 1 0 resetb $end
$var wire 1 ' rx $end
$var wire 1 ( tx $end
$var wire 1 " host_dor $end
$var wire 1 # host_dir $end
$var reg 2 D din_q [1:0] $end
$var reg 32 E par2ser_q [31:0] $end
$var reg 1 F rx_ack_req_q $end
$var reg 5 G rx_count_q [4:0] $end
$var reg 1 H rx_ready_q $end
$var reg 2 I rx_state_q [1:0] $end
$var reg 32 J ser2par_q [31:0] $end
$var reg 1 K tx_ack_rcvd_q $end
$var reg 5 L tx_count_q [4:0] $end
$var reg 1 M tx_r $end
$var reg 1 N tx_ready_q $end
$var reg 3 O tx_state_q [2:0] $end
$upscope $end
$scope task transmitAB $end
$var reg 32 P data [31:0] $end
$upscope $end
$scope task transmitBA $end
$var reg 32 Q data [31:0] $end
$upscope $end
$upscope $end
$enddefinitions $end
#0
$dumpvars
bx Q
bx P
b0 O
0N
0M
b0 L
0K
b0 J
b0 I
1H
b0 G
0F
b0 E
b0 D
b0 C
bx B
b0 A
b0 @
0?
0>
b0 =
0<
b0 ;
b0 :
19
b0 8
07
b0 6
b0 5
b0 4
bx 3
b0 2
01
00
0/
0.
bx -
0,
0+
bx *
0)
0(
0'
1&
0%
b0 $
1#
0"
b0 !
$end
#100
1)
#200
0)
#300
1)
#400
0)
#500
1)
#600
0)
#700
1)
#800
0)
#900
1)
#1000
0)
#1100
10
1)
#1200
0)
#1300
1)
#1400
0)
#1500
1)
#1600
0)
#1700
1)
#1800
0)
#1900
1)
#2000
0)
#2100
0&
1?
1,
1)
b1001000110100010101100111 *
b1001000110100010101100111 3
b1001000110100010101100111 P
#2200
b1001000110100010101100111 6
0)
#2300
1'
1>
b100 @
0,
1)
#2400
b1 A
b1 D
0)
#2500
b101 @
1)
#2600
b11 A
b11 D
0)
#2700
0'
0>
b10 @
b10 I
1)
#2800
b10010001101000101011001110 6
b10 A
b10 D
0)
#2900
b1 G
b1 =
1)
#3000
b0 A
b0 D
b100100011010001010110011100 6
0)
#3100
b10 =
b10 G
1)
#3200
b1001000110100010101100111000 6
0)
#3300
b11 G
b11 =
1)
#3400
b10010001101000101011001110000 6
0)
#3500
b100 =
b100 G
1)
#3600
b100100011010001010110011100000 6
0)
#3700
b101 G
b101 =
1)
#3800
b1001000110100010101100111000000 6
0)
#3900
b110 =
b110 G
1)
#4000
1'
1>
b10010001101000101011001110000000 6
0)
#4100
b111 G
b111 =
1)
#4200
0'
0>
b1 A
b1 D
b1 !
b1 C
b1 J
b100011010001010110011100000000 6
0)
#4300
b1000 =
b1000 G
1)
#4400
b1000110100010101100111000000000 6
b10 A
b10 D
b10 !
b10 C
b10 J
0)
#4500
b1001 G
b1001 =
1)
#4600
1'
1>
b0 A
b0 D
b100 !
b100 C
b100 J
b10001101000101011001110000000000 6
0)
#4700
b1010 =
b1010 G
1)
#4800
0'
0>
b11010001010110011100000000000 6
b1 A
b1 D
b1001 !
b1001 C
b1001 J
0)
#4900
b1011 G
b1011 =
1)
#5000
b10 A
b10 D
b10010 !
b10010 C
b10010 J
b110100010101100111000000000000 6
0)
#5100
b1100 =
b1100 G
1)
#5200
b1101000101011001110000000000000 6
b0 A
b0 D
b100100 !
b100100 C
b100100 J
0)
#5300
b1101 G
b1101 =
1)
#5400
1'
1>
b1001000 !
b1001000 C
b1001000 J
b11010001010110011100000000000000 6
0)
#5500
b1110 =
b1110 G
1)
#5600
b10100010101100111000000000000000 6
b1 A
b1 D
b10010001 !
b10010001 C
b10010001 J
0)
#5700
b1111 G
b1111 =
1)
#5800
0'
0>
b11 A
b11 D
b100100011 !
b100100011 C
b100100011 J
b1000101011001110000000000000000 6
0)
#5900
b10000 =
b10000 G
1)
#6000
1'
1>
b10001010110011100000000000000000 6
b10 A
b10 D
b1001000110 !
b1001000110 C
b1001000110 J
0)
#6100
b10001 G
b10001 =
1)
#6200
0'
0>
b1 A
b1 D
b10010001101 !
b10010001101 C
b10010001101 J
b10101100111000000000000000000 6
0)
#6300
b10010 =
b10010 G
1)
#6400
b101011001110000000000000000000 6
b10 A
b10 D
b100100011010 !
b100100011010 C
b100100011010 J
0)
#6500
b10011 G
b10011 =
1)
#6600
b0 A
b0 D
b1001000110100 !
b1001000110100 C
b1001000110100 J
b1010110011100000000000000000000 6
0)
#6700
b10100 =
b10100 G
1)
#6800
1'
1>
b10101100111000000000000000000000 6
b10010001101000 !
b10010001101000 C
b10010001101000 J
0)
#6900
b10101 G
b10101 =
1)
#7000
0'
0>
b1 A
b1 D
b100100011010001 !
b100100011010001 C
b100100011010001 J
b1011001110000000000000000000000 6
0)
#7100
b10110 =
b10110 G
1)
#7200
1'
1>
b10110011100000000000000000000000 6
b10 A
b10 D
b1001000110100010 !
b1001000110100010 C
b1001000110100010 J
0)
#7300
b10111 G
b10111 =
1)
#7400
0'
0>
b1 A
b1 D
b10010001101000101 !
b10010001101000101 C
b10010001101000101 J
b1100111000000000000000000000000 6
0)
#7500
b11000 =
b11000 G
1)
#7600
1'
1>
b11001110000000000000000000000000 6
b10 A
b10 D
b100100011010001010 !
b100100011010001010 C
b100100011010001010 J
0)
#7700
b11001 G
b11001 =
1)
#7800
b1 A
b1 D
b1001000110100010101 !
b1001000110100010101 C
b1001000110100010101 J
b10011100000000000000000000000000 6
0)
#7900
b11010 =
b11010 G
1)
#8000
0'
0>
b111000000000000000000000000000 6
b11 A
b11 D
b10010001101000101011 !
b10010001101000101011 C
b10010001101000101011 J
0)
#8100
b11011 G
b11011 =
1)
#8200
b10 A
b10 D
b100100011010001010110 !
b100100011010001010110 C
b100100011010001010110 J
b1110000000000000000000000000000 6
0)
#8300
b11100 =
b11100 G
1)
#8400
1'
1>
b11100000000000000000000000000000 6
b0 A
b0 D
b1001000110100010101100 !
b1001000110100010101100 C
b1001000110100010101100 J
0)
#8500
b11101 G
b11101 =
1)
#8600
b1 A
b1 D
b10010001101000101011001 !
b10010001101000101011001 C
b10010001101000101011001 J
b11000000000000000000000000000000 6
0)
#8700
b11110 =
b11110 G
1)
#8800
b10000000000000000000000000000000 6
b11 A
b11 D
b100100011010001010110011 !
b100100011010001010110011 C
b100100011010001010110011 J
0)
#8900
b11111 G
b11111 =
1)
#9000
0'
0>
b1001000110100010101100111 !
b1001000110100010101100111 C
b1001000110100010101100111 J
b0 6
0)
#9100
b11 @
b0 =
b11 I
b0 G
1)
#9200
b10 A
b10 D
0)
#9300
1"
0H
1F
b1 I
1)
#9400
b0 A
b0 D
0)
#9500
1(
1M
b110 O
b0 I
1)
#9600
b1 2
b1 5
0)
#9700
0(
0M
0"
1H
b111 O
1.
1)
#9800
b10 2
b10 5
0)
#9900
1<
b0 O
0F
b10001001101010111100110111101111 *
b10001001101010111100110111101111 3
b10001001101010111100110111101111 P
0.
1)
#10000
b0 2
b0 5
0)
#10100
b1 @
1)
#10200
0)
#10300
b0 @
1&
0?
1)
#10400
0)
#10500
1)
#10600
0)
#10700
0&
1?
1,
1)
#10800
b10001001101010111100110111101111 6
0)
#10900
1'
1>
b100 @
0,
1)
#11000
b1 A
b1 D
0)
#11100
b101 @
0<
1)
#11200
b11 A
b11 D
0)
#11300
b10 I
b10 @
1)
#11400
0'
0>
b10010001101000101011001111 !
b10010001101000101011001111 C
b10010001101000101011001111 J
b10011010101111001101111011110 6
0)
#11500
b1 =
b1 G
1)
#11600
b100110101011110011011110111100 6
b10 A
b10 D
b100100011010001010110011110 !
b100100011010001010110011110 C
b100100011010001010110011110 J
0)
#11700
b10 G
b10 =
1)
#11800
b0 A
b0 D
b1001000110100010101100111100 !
b1001000110100010101100111100 C
b1001000110100010101100111100 J
b1001101010111100110111101111000 6
0)
#11900
b11 =
b11 G
1)
#12000
1'
1>
b10011010101111001101111011110000 6
b10010001101000101011001111000 !
b10010001101000101011001111000 C
b10010001101000101011001111000 J
0)
#12100
b100 G
b100 =
1)
#12200
0'
0>
b1 A
b1 D
b100100011010001010110011110001 !
b100100011010001010110011110001 C
b100100011010001010110011110001 J
b110101011110011011110111100000 6
0)
#12300
b101 =
b101 G
1)
#12400
b1101010111100110111101111000000 6
b10 A
b10 D
b1001000110100010101100111100010 !
b1001000110100010101100111100010 C
b1001000110100010101100111100010 J
0)
#12500
b110 G
b110 =
1)
#12600
1'
1>
b0 A
b0 D
b10010001101000101011001111000100 !
b10010001101000101011001111000100 C
b10010001101000101011001111000100 J
b11010101111001101111011110000000 6
0)
#12700
b111 =
b111 G
1)
#12800
b10101011110011011110111100000000 6
b1 A
b1 D
b100011010001010110011110001001 !
b100011010001010110011110001001 C
b100011010001010110011110001001 J
0)
#12900
b1000 G
b1000 =
1)
#13000
0'
0>
b11 A
b11 D
b1000110100010101100111100010011 !
b1000110100010101100111100010011 C
b1000110100010101100111100010011 J
b1010111100110111101111000000000 6
0)
#13100
b1001 =
b1001 G
1)
#13200
1'
1>
b10101111001101111011110000000000 6
b10 A
b10 D
b10001101000101011001111000100110 !
b10001101000101011001111000100110 C
b10001101000101011001111000100110 J
0)
#13300
b1010 G
b1010 =
1)
#13400
0'
0>
b1 A
b1 D
b11010001010110011110001001101 !
b11010001010110011110001001101 C
b11010001010110011110001001101 J
b1011110011011110111100000000000 6
0)
#13500
b1011 =
b1011 G
1)
#13600
1'
1>
b10111100110111101111000000000000 6
b10 A
b10 D
b110100010101100111100010011010 !
b110100010101100111100010011010 C
b110100010101100111100010011010 J
0)
#13700
b1100 G
b1100 =
1)
#13800
0'
0>
b1 A
b1 D
b1101000101011001111000100110101 !
b1101000101011001111000100110101 C
b1101000101011001111000100110101 J
b1111001101111011110000000000000 6
0)
#13900
b1101 =
b1101 G
1)
#14000
1'
1>
b11110011011110111100000000000000 6
b10 A
b10 D
b11010001010110011110001001101010 !
b11010001010110011110001001101010 C
b11010001010110011110001001101010 J
0)
#14100
b1110 G
b1110 =
1)
#14200
b1 A
b1 D
b10100010101100111100010011010101 !
b10100010101100111100010011010101 C
b10100010101100111100010011010101 J
b11100110111101111000000000000000 6
0)
#14300
b1111 =
b1111 G
1)
#14400
b11001101111011110000000000000000 6
b11 A
b11 D
b1000101011001111000100110101011 !
b1000101011001111000100110101011 C
b1000101011001111000100110101011 J
0)
#14500
b10000 G
b10000 =
1)
#14600
b10001010110011110001001101010111 !
b10001010110011110001001101010111 C
b10001010110011110001001101010111 J
b10011011110111100000000000000000 6
0)
#14700
b10001 =
b10001 G
1)
#14800
0'
0>
b110111101111000000000000000000 6
b10101100111100010011010101111 !
b10101100111100010011010101111 C
b10101100111100010011010101111 J
0)
#14900
b10010 G
b10010 =
1)
#15000
b10 A
b10 D
b101011001111000100110101011110 !
b101011001111000100110101011110 C
b101011001111000100110101011110 J
b1101111011110000000000000000000 6
0)
#15100
b10011 =
b10011 G
1)
#15200
1'
1>
b11011110111100000000000000000000 6
b0 A
b0 D
b1010110011110001001101010111100 !
b1010110011110001001101010111100 C
b1010110011110001001101010111100 J
0)
#15300
b10100 G
b10100 =
1)
#15400
b1 A
b1 D
b10101100111100010011010101111001 !
b10101100111100010011010101111001 C
b10101100111100010011010101111001 J
b10111101111000000000000000000000 6
0)
#15500
b10101 =
b10101 G
1)
#15600
0'
0>
b1111011110000000000000000000000 6
b11 A
b11 D
b1011001111000100110101011110011 !
b1011001111000100110101011110011 C
b1011001111000100110101011110011 J
0)
#15700
b10110 G
b10110 =
1)
#15800
1'
1>
b10 A
b10 D
b10110011110001001101010111100110 !
b10110011110001001101010111100110 C
b10110011110001001101010111100110 J
b11110111100000000000000000000000 6
0)
#15900
b10111 =
b10111 G
1)
#16000
b11101111000000000000000000000000 6
b1 A
b1 D
b1100111100010011010101111001101 !
b1100111100010011010101111001101 C
b1100111100010011010101111001101 J
0)
#16100
b11000 G
b11000 =
1)
#16200
b11 A
b11 D
b11001111000100110101011110011011 !
b11001111000100110101011110011011 C
b11001111000100110101011110011011 J
b11011110000000000000000000000000 6
0)
#16300
b11001 =
b11001 G
1)
#16400
b10111100000000000000000000000000 6
b10011110001001101010111100110111 !
b10011110001001101010111100110111 C
b10011110001001101010111100110111 J
0)
#16500
b11010 G
b11010 =
1)
#16600
0'
0>
b111100010011010101111001101111 !
b111100010011010101111001101111 C
b111100010011010101111001101111 J
b1111000000000000000000000000000 6
0)
#16700
b11011 =
b11011 G
1)
#16800
1'
1>
b11110000000000000000000000000000 6
b10 A
b10 D
b1111000100110101011110011011110 !
b1111000100110101011110011011110 C
b1111000100110101011110011011110 J
0)
#16900
b11100 G
b11100 =
1)
#17000
b1 A
b1 D
b11110001001101010111100110111101 !
b11110001001101010111100110111101 C
b11110001001101010111100110111101 J
b11100000000000000000000000000000 6
0)
#17100
b11101 =
b11101 G
1)
#17200
b11000000000000000000000000000000 6
b11 A
b11 D
b11100010011010101111001101111011 !
b11100010011010101111001101111011 C
b11100010011010101111001101111011 J
0)
#17300
b11110 G
b11110 =
1)
#17400
b11000100110101011110011011110111 !
b11000100110101011110011011110111 C
b11000100110101011110011011110111 J
b10000000000000000000000000000000 6
0)
#17500
b11111 =
b11111 G
1)
#17600
0'
0>
b0 6
b10001001101010111100110111101111 !
b10001001101010111100110111101111 C
b10001001101010111100110111101111 J
0)
#17700
b0 G
b11 I
b0 =
b11 @
1)
#17800
b10 A
b10 D
0)
#17900
b1 I
1F
1"
0H
1)
#18000
b0 A
b0 D
0)
#18100
1(
1M
b0 I
b110 O
1)
#18200
b1 2
b1 5
0)
#18300
0(
0M
b111 O
0"
1H
1.
1)
#18400
b10 2
b10 5
0)
#18500
0F
b0 O
1<
b100010010001000110011 *
b100010010001000110011 3
b100010010001000110011 P
0.
1)
#18600
b0 2
b0 5
0)
#18700
b1 @
1)
#18800
0)
#18900
1&
0?
b0 @
1)
#19000
0)
#19100
1)
#19200
0)
#19300
0&
1?
1,
1)
#19400
b100010010001000110011 6
0)
#19500
1'
1>
b100 @
0,
1)
#19600
b1 A
b1 D
0)
#19700
0<
b101 @
1)
#19800
b11 A
b11 D
0)
#19900
0'
0>
b10 @
b10 I
1)
#20000
b1000100100010001100110 6
b10 A
b10 D
b10011010101111001101111011110 !
b10011010101111001101111011110 C
b10011010101111001101111011110 J
0)
#20100
b1 G
b1 =
1)
#20200
b0 A
b0 D
b100110101011110011011110111100 !
b100110101011110011011110111100 C
b100110101011110011011110111100 J
b10001001000100011001100 6
0)
#20300
b10 =
b10 G
1)
#20400
b100010010001000110011000 6
b1001101010111100110111101111000 !
b1001101010111100110111101111000 C
b1001101010111100110111101111000 J
0)
#20500
b11 G
b11 =
1)
#20600
b10011010101111001101111011110000 !
b10011010101111001101111011110000 C
b10011010101111001101111011110000 J
b1000100100010001100110000 6
0)
#20700
b100 =
b100 G
1)
#20800
b10001001000100011001100000 6
b110101011110011011110111100000 !
b110101011110011011110111100000 C
b110101011110011011110111100000 J
0)
#20900
b101 G
b101 =
1)
#21000
b1101010111100110111101111000000 !
b1101010111100110111101111000000 C
b1101010111100110111101111000000 J
b100010010001000110011000000 6
0)
#21100
b110 =
b110 G
1)
#21200
b1000100100010001100110000000 6
b11010101111001101111011110000000 !
b11010101111001101111011110000000 C
b11010101111001101111011110000000 J
0)
#21300
b111 G
b111 =
1)
#21400
b10101011110011011110111100000000 !
b10101011110011011110111100000000 C
b10101011110011011110111100000000 J
b10001001000100011001100000000 6
0)
#21500
b1000 =
b1000 G
1)
#21600
b100010010001000110011000000000 6
b1010111100110111101111000000000 !
b1010111100110111101111000000000 C
b1010111100110111101111000000000 J
0)
#21700
b1001 G
b1001 =
1)
#21800
b10101111001101111011110000000000 !
b10101111001101111011110000000000 C
b10101111001101111011110000000000 J
b1000100100010001100110000000000 6
0)
#21900
b1010 =
b1010 G
1)
#22000
1'
1>
b10001001000100011001100000000000 6
b1011110011011110111100000000000 !
b1011110011011110111100000000000 C
b1011110011011110111100000000000 J
0)
#22100
b1011 G
b1011 =
1)
#22200
0'
0>
b1 A
b1 D
b10111100110111101111000000000001 !
b10111100110111101111000000000001 C
b10111100110111101111000000000001 J
b10010001000110011000000000000 6
0)
#22300
b1100 =
b1100 G
1)
#22400
b100100010001100110000000000000 6
b10 A
b10 D
b1111001101111011110000000000010 !
b1111001101111011110000000000010 C
b1111001101111011110000000000010 J
0)
#22500
b1101 G
b1101 =
1)
#22600
b0 A
b0 D
b11110011011110111100000000000100 !
b11110011011110111100000000000100 C
b11110011011110111100000000000100 J
b1001000100011001100000000000000 6
0)
#22700
b1110 =
b1110 G
1)
#22800
1'
1>
b10010001000110011000000000000000 6
b11100110111101111000000000001000 !
b11100110111101111000000000001000 C
b11100110111101111000000000001000 J
0)
#22900
b1111 G
b1111 =
1)
#23000
0'
0>
b1 A
b1 D
b11001101111011110000000000010001 !
b11001101111011110000000000010001 C
b11001101111011110000000000010001 J
b100010001100110000000000000000 6
0)
#23100
b10000 =
b10000 G
1)
#23200
b1000100011001100000000000000000 6
b10 A
b10 D
b10011011110111100000000000100010 !
b10011011110111100000000000100010 C
b10011011110111100000000000100010 J
0)
#23300
b10001 G
b10001 =
1)
#23400
1'
1>
b0 A
b0 D
b110111101111000000000001000100 !
b110111101111000000000001000100 C
b110111101111000000000001000100 J
b10001000110011000000000000000000 6
0)
#23500
b10010 =
b10010 G
1)
#23600
0'
0>
b10001100110000000000000000000 6
b1 A
b1 D
b1101111011110000000000010001001 !
b1101111011110000000000010001001 C
b1101111011110000000000010001001 J
0)
#23700
b10011 G
b10011 =
1)
#23800
b10 A
b10 D
b11011110111100000000000100010010 !
b11011110111100000000000100010010 C
b11011110111100000000000100010010 J
b100011001100000000000000000000 6
0)
#23900
b10100 =
b10100 G
1)
#24000
b1000110011000000000000000000000 6
b0 A
b0 D
b10111101111000000000001000100100 !
b10111101111000000000001000100100 C
b10111101111000000000001000100100 J
0)
#24100
b10101 G
b10101 =
1)
#24200
1'
1>
b1111011110000000000010001001000 !
b1111011110000000000010001001000 C
b1111011110000000000010001001000 J
b10001100110000000000000000000000 6
0)
#24300
b10110 =
b10110 G
1)
#24400
0'
0>
b11001100000000000000000000000 6
b1 A
b1 D
b11110111100000000000100010010001 !
b11110111100000000000100010010001 C
b11110111100000000000100010010001 J
0)
#24500
b10111 G
b10111 =
1)
#24600
b10 A
b10 D
b11101111000000000001000100100010 !
b11101111000000000001000100100010 C
b11101111000000000001000100100010 J
b110011000000000000000000000000 6
0)
#24700
b11000 =
b11000 G
1)
#24800
b1100110000000000000000000000000 6
b0 A
b0 D
b11011110000000000010001001000100 !
b11011110000000000010001001000100 C
b11011110000000000010001001000100 J
0)
#24900
b11001 G
b11001 =
1)
#25000
1'
1>
b10111100000000000100010010001000 !
b10111100000000000100010010001000 C
b10111100000000000100010010001000 J
b11001100000000000000000000000000 6
0)
#25100
b11010 =
b11010 G
1)
#25200
b10011000000000000000000000000000 6
b1 A
b1 D
b1111000000000001000100100010001 !
b1111000000000001000100100010001 C
b1111000000000001000100100010001 J
0)
#25300
b11011 G
b11011 =
1)
#25400
0'
0>
b11 A
b11 D
b11110000000000010001001000100011 !
b11110000000000010001001000100011 C
b11110000000000010001001000100011 J
b110000000000000000000000000000 6
0)
#25500
b11100 =
b11100 G
1)
#25600
b1100000000000000000000000000000 6
b10 A
b10 D
b11100000000000100010010001000110 !
b11100000000000100010010001000110 C
b11100000000000100010010001000110 J
0)
#25700
b11101 G
b11101 =
1)
#25800
1'
1>
b0 A
b0 D
b11000000000001000100100010001100 !
b11000000000001000100100010001100 C
b11000000000001000100100010001100 J
b11000000000000000000000000000000 6
0)
#25900
b11110 =
b11110 G
1)
#26000
b10000000000000000000000000000000 6
b1 A
b1 D
b10000000000010001001000100011001 !
b10000000000010001001000100011001 C
b10000000000010001001000100011001 J
0)
#26100
b11111 G
b11111 =
1)
#26200
0'
0>
b11 A
b11 D
b100010010001000110011 !
b100010010001000110011 C
b100010010001000110011 J
b0 6
0)
#26300
b11 @
b0 =
b11 I
b0 G
1)
#26400
b10 A
b10 D
0)
#26500
1"
0H
1F
b1 I
1)
#26600
b0 A
b0 D
0)
#26700
1(
1M
b110 O
b0 I
1)
#26800
b1 2
b1 5
0)
#26900
0(
0M
0"
1H
b111 O
1.
1)
#27000
b10 2
b10 5
0)
#27100
1<
b0 O
0F
b1000100010101010110011001110111 *
b1000100010101010110011001110111 3
b1000100010101010110011001110111 P
0.
1)
#27200
b0 2
b0 5
0)
#27300
b1 @
1)
#27400
0)
#27500
b0 @
1&
0?
1)
#27600
0)
#27700
1)
#27800
0)
#27900
0&
1?
1,
1)
#28000
b1000100010101010110011001110111 6
0)
#28100
1'
1>
b100 @
0,
1)
#28200
b1 A
b1 D
0)
#28300
b101 @
0<
1)
#28400
b11 A
b11 D
0)
#28500
0'
0>
b10 I
b10 @
1)
#28600
1'
1>
b10 A
b10 D
b1000100100010001100110 !
b1000100100010001100110 C
b1000100100010001100110 J
b10001000101010101100110011101110 6
0)
#28700
b1 =
b1 G
1)
#28800
0'
0>
b10001010101011001100111011100 6
b1 A
b1 D
b10001001000100011001101 !
b10001001000100011001101 C
b10001001000100011001101 J
0)
#28900
b10 G
b10 =
1)
#29000
b10 A
b10 D
b100010010001000110011010 !
b100010010001000110011010 C
b100010010001000110011010 J
b100010101010110011001110111000 6
0)
#29100
b11 =
b11 G
1)
#29200
b1000101010101100110011101110000 6
b0 A
b0 D
b1000100100010001100110100 !
b1000100100010001100110100 C
b1000100100010001100110100 J
0)
#29300
b100 G
b100 =
1)
#29400
1'
1>
b10001001000100011001101000 !
b10001001000100011001101000 C
b10001001000100011001101000 J
b10001010101011001100111011100000 6
0)
#29500
b101 =
b101 G
1)
#29600
0'
0>
b10101010110011001110111000000 6
b1 A
b1 D
b100010010001000110011010001 !
b100010010001000110011010001 C
b100010010001000110011010001 J
0)
#29700
b110 G
b110 =
1)
#29800
b10 A
b10 D
b1000100100010001100110100010 !
b1000100100010001100110100010 C
b1000100100010001100110100010 J
b101010101100110011101110000000 6
0)
#29900
b111 =
b111 G
1)
#30000
b1010101011001100111011100000000 6
b0 A
b0 D
b10001001000100011001101000100 !
b10001001000100011001101000100 C
b10001001000100011001101000100 J
0)
#30100
b1000 G
b1000 =
1)
#30200
1'
1>
b100010010001000110011010001000 !
b100010010001000110011010001000 C
b100010010001000110011010001000 J
b10101010110011001110111000000000 6
0)
#30300
b1001 =
b1001 G
1)
#30400
0'
0>
b1010101100110011101110000000000 6
b1 A
b1 D
b1000100100010001100110100010001 !
b1000100100010001100110100010001 C
b1000100100010001100110100010001 J
0)
#30500
b1010 G
b1010 =
1)
#30600
1'
1>
b10 A
b10 D
b10001001000100011001101000100010 !
b10001001000100011001101000100010 C
b10001001000100011001101000100010 J
b10101011001100111011100000000000 6
0)
#30700
b1011 =
b1011 G
1)
#30800
0'
0>
b1010110011001110111000000000000 6
b1 A
b1 D
b10010001000110011010001000101 !
b10010001000110011010001000101 C
b10010001000110011010001000101 J
0)
#30900
b1100 G
b1100 =
1)
#31000
1'
1>
b10 A
b10 D
b100100010001100110100010001010 !
b100100010001100110100010001010 C
b100100010001100110100010001010 J
b10101100110011101110000000000000 6
0)
#31100
b1101 =
b1101 G
1)
#31200
0'
0>
b1011001100111011100000000000000 6
b1 A
b1 D
b1001000100011001101000100010101 !
b1001000100011001101000100010101 C
b1001000100011001101000100010101 J
0)
#31300
b1110 G
b1110 =
1)
#31400
1'
1>
b10 A
b10 D
b10010001000110011010001000101010 !
b10010001000110011010001000101010 C
b10010001000110011010001000101010 J
b10110011001110111000000000000000 6
0)
#31500
b1111 =
b1111 G
1)
#31600
0'
0>
b1100110011101110000000000000000 6
b1 A
b1 D
b100010001100110100010001010101 !
b100010001100110100010001010101 C
b100010001100110100010001010101 J
0)
#31700
b10000 G
b10000 =
1)
#31800
1'
1>
b10 A
b10 D
b1000100011001101000100010101010 !
b1000100011001101000100010101010 C
b1000100011001101000100010101010 J
b11001100111011100000000000000000 6
0)
#31900
b10001 =
b10001 G
1)
#32000
b10011001110111000000000000000000 6
b1 A
b1 D
b10001000110011010001000101010101 !
b10001000110011010001000101010101 C
b10001000110011010001000101010101 J
0)
#32100
b10010 G
b10010 =
1)
#32200
0'
0>
b11 A
b11 D
b10001100110100010001010101011 !
b10001100110100010001010101011 C
b10001100110100010001010101011 J
b110011101110000000000000000000 6
0)
#32300
b10011 =
b10011 G
1)
#32400
b1100111011100000000000000000000 6
b10 A
b10 D
b100011001101000100010101010110 !
b100011001101000100010101010110 C
b100011001101000100010101010110 J
0)
#32500
b10100 G
b10100 =
1)
#32600
1'
1>
b0 A
b0 D
b1000110011010001000101010101100 !
b1000110011010001000101010101100 C
b1000110011010001000101010101100 J
b11001110111000000000000000000000 6
0)
#32700
b10101 =
b10101 G
1)
#32800
b10011101110000000000000000000000 6
b1 A
b1 D
b10001100110100010001010101011001 !
b10001100110100010001010101011001 C
b10001100110100010001010101011001 J
0)
#32900
b10110 G
b10110 =
1)
#33000
0'
0>
b11 A
b11 D
b11001101000100010101010110011 !
b11001101000100010101010110011 C
b11001101000100010101010110011 J
b111011100000000000000000000000 6
0)
#33100
b10111 =
b10111 G
1)
#33200
b1110111000000000000000000000000 6
b10 A
b10 D
b110011010001000101010101100110 !
b110011010001000101010101100110 C
b110011010001000101010101100110 J
0)
#33300
b11000 G
b11000 =
1)
#33400
1'
1>
b0 A
b0 D
b1100110100010001010101011001100 !
b1100110100010001010101011001100 C
b1100110100010001010101011001100 J
b11101110000000000000000000000000 6
0)
#33500
b11001 =
b11001 G
1)
#33600
b11011100000000000000000000000000 6
b1 A
b1 D
b11001101000100010101010110011001 !
b11001101000100010101010110011001 C
b11001101000100010101010110011001 J
0)
#33700
b11010 G
b11010 =
1)
#33800
b11 A
b11 D
b10011010001000101010101100110011 !
b10011010001000101010101100110011 C
b10011010001000101010101100110011 J
b10111000000000000000000000000000 6
0)
#33900
b11011 =
b11011 G
1)
#34000
0'
0>
b1110000000000000000000000000000 6
b110100010001010101011001100111 !
b110100010001010101011001100111 C
b110100010001010101011001100111 J
0)
#34100
b11100 G
b11100 =
1)
#34200
1'
1>
b10 A
b10 D
b1101000100010101010110011001110 !
b1101000100010101010110011001110 C
b1101000100010101010110011001110 J
b11100000000000000000000000000000 6
0)
#34300
b11101 =
b11101 G
1)
#34400
b11000000000000000000000000000000 6
b1 A
b1 D
b11010001000101010101100110011101 !
b11010001000101010101100110011101 C
b11010001000101010101100110011101 J
0)
#34500
b11110 G
b11110 =
1)
#34600
b11 A
b11 D
b10100010001010101011001100111011 !
b10100010001010101011001100111011 C
b10100010001010101011001100111011 J
b10000000000000000000000000000000 6
0)
#34700
b11111 =
b11111 G
1)
#34800
0'
0>
b0 6
b1000100010101010110011001110111 !
b1000100010101010110011001110111 C
b1000100010101010110011001110111 J
0)
#34900
b0 G
b11 I
b0 =
b11 @
1)
#35000
b10 A
b10 D
0)
#35100
b1 I
1F
1"
0H
1)
#35200
b0 A
b0 D
0)
#35300
1(
1M
b0 I
b110 O
1)
#35400
b1 2
b1 5
0)
#35500
0(
0M
b111 O
0"
1H
1.
1)
#35600
b10 2
b10 5
0)
#35700
0F
b0 O
1<
b1001000110100010101100111 -
b1001000110100010101100111 B
b1001000110100010101100111 Q
0.
1)
#35800
b0 2
b0 5
0)
#35900
b1 @
0#
1N
1/
1)
#36000
b1001000110100010101100111 E
0)
#36100
1(
1M
b100 O
1&
0?
b0 @
0/
1)
#36200
b1 2
b1 5
0)
#36300
b101 O
1)
#36400
b11 2
b11 5
0)
#36500
0(
0M
b10 O
b10 :
1)
#36600
b10010001101000101011001110 E
b10 2
b10 5
0)
#36700
b1 8
b1 L
1)
#36800
b0 2
b0 5
b100100011010001010110011100 E
0)
#36900
b10 L
b10 8
1)
#37000
b1001000110100010101100111000 E
0)
#37100
b11 8
b11 L
1)
#37200
b10010001101000101011001110000 E
0)
#37300
b100 L
b100 8
1)
#37400
b100100011010001010110011100000 E
0)
#37500
b101 8
b101 L
1)
#37600
b1001000110100010101100111000000 E
0)
#37700
b110 L
b110 8
1)
#37800
1(
1M
b10010001101000101011001110000000 E
0)
#37900
b111 8
b111 L
1)
#38000
0(
0M
b1 2
b1 5
b1 $
b1 4
b1 ;
b100011010001010110011100000000 E
0)
#38100
b1000 L
b1000 8
1)
#38200
b1000110100010101100111000000000 E
b10 2
b10 5
b10 $
b10 4
b10 ;
0)
#38300
b1001 8
b1001 L
1)
#38400
1(
1M
b0 2
b0 5
b100 $
b100 4
b100 ;
b10001101000101011001110000000000 E
0)
#38500
b1010 L
b1010 8
1)
#38600
0(
0M
b11010001010110011100000000000 E
b1 2
b1 5
b1001 $
b1001 4
b1001 ;
0)
#38700
b1011 8
b1011 L
1)
#38800
b10 2
b10 5
b10010 $
b10010 4
b10010 ;
b110100010101100111000000000000 E
0)
#38900
b1100 L
b1100 8
1)
#39000
b1101000101011001110000000000000 E
b0 2
b0 5
b100100 $
b100100 4
b100100 ;
0)
#39100
b1101 8
b1101 L
1)
#39200
1(
1M
b1001000 $
b1001000 4
b1001000 ;
b11010001010110011100000000000000 E
0)
#39300
b1110 L
b1110 8
1)
#39400
b10100010101100111000000000000000 E
b1 2
b1 5
b10010001 $
b10010001 4
b10010001 ;
0)
#39500
b1111 8
b1111 L
1)
#39600
0(
0M
b11 2
b11 5
b100100011 $
b100100011 4
b100100011 ;
b1000101011001110000000000000000 E
0)
#39700
b10000 L
b10000 8
1)
#39800
1(
1M
b10001010110011100000000000000000 E
b10 2
b10 5
b1001000110 $
b1001000110 4
b1001000110 ;
0)
#39900
b10001 8
b10001 L
1)
#40000
0(
0M
b1 2
b1 5
b10010001101 $
b10010001101 4
b10010001101 ;
b10101100111000000000000000000 E
0)
#40100
b10010 L
b10010 8
1)
#40200
b101011001110000000000000000000 E
b10 2
b10 5
b100100011010 $
b100100011010 4
b100100011010 ;
0)
#40300
b10011 8
b10011 L
1)
#40400
b0 2
b0 5
b1001000110100 $
b1001000110100 4
b1001000110100 ;
b1010110011100000000000000000000 E
0)
#40500
b10100 L
b10100 8
1)
#40600
1(
1M
b10101100111000000000000000000000 E
b10010001101000 $
b10010001101000 4
b10010001101000 ;
0)
#40700
b10101 8
b10101 L
1)
#40800
0(
0M
b1 2
b1 5
b100100011010001 $
b100100011010001 4
b100100011010001 ;
b1011001110000000000000000000000 E
0)
#40900
b10110 L
b10110 8
1)
#41000
1(
1M
b10110011100000000000000000000000 E
b10 2
b10 5
b1001000110100010 $
b1001000110100010 4
b1001000110100010 ;
0)
#41100
b10111 8
b10111 L
1)
#41200
0(
0M
b1 2
b1 5
b10010001101000101 $
b10010001101000101 4
b10010001101000101 ;
b1100111000000000000000000000000 E
0)
#41300
b11000 L
b11000 8
1)
#41400
1(
1M
b11001110000000000000000000000000 E
b10 2
b10 5
b100100011010001010 $
b100100011010001010 4
b100100011010001010 ;
0)
#41500
b11001 8
b11001 L
1)
#41600
b1 2
b1 5
b1001000110100010101 $
b1001000110100010101 4
b1001000110100010101 ;
b10011100000000000000000000000000 E
0)
#41700
b11010 L
b11010 8
1)
#41800
0(
0M
b111000000000000000000000000000 E
b11 2
b11 5
b10010001101000101011 $
b10010001101000101011 4
b10010001101000101011 ;
0)
#41900
b11011 8
b11011 L
1)
#42000
b10 2
b10 5
b100100011010001010110 $
b100100011010001010110 4
b100100011010001010110 ;
b1110000000000000000000000000000 E
0)
#42100
b11100 L
b11100 8
1)
#42200
1(
1M
b11100000000000000000000000000000 E
b0 2
b0 5
b1001000110100010101100 $
b1001000110100010101100 4
b1001000110100010101100 ;
0)
#42300
b11101 8
b11101 L
1)
#42400
b1 2
b1 5
b10010001101000101011001 $
b10010001101000101011001 4
b10010001101000101011001 ;
b11000000000000000000000000000000 E
0)
#42500
b11110 L
b11110 8
1)
#42600
b10000000000000000000000000000000 E
b11 2
b11 5
b100100011010001010110011 $
b100100011010001010110011 4
b100100011010001010110011 ;
0)
#42700
b11111 8
b11111 L
1)
#42800
0(
0M
b1001000110100010101100111 $
b1001000110100010101100111 4
b1001000110100010101100111 ;
b0 E
0)
#42900
b0 L
b11 O
b0 8
b11 :
1)
#43000
b10 2
b10 5
0)
#43100
b1 :
17
1%
09
1)
#43200
b0 2
b0 5
0)
#43300
1'
1>
b0 :
b110 @
1)
#43400
b1 A
b1 D
0)
#43500
0'
0>
b111 @
0%
19
1+
1)
#43600
b10 A
b10 D
0)
#43700
1K
07
b0 @
b10001001101010111100110111101111 -
b10001001101010111100110111101111 B
b10001001101010111100110111101111 Q
0+
1)
#43800
b0 A
b0 D
0)
#43900
b1 O
1)
#44000
0)
#44100
1#
0N
b0 O
1)
#44200
0)
#44300
1)
#44400
0)
#44500
0#
1N
1/
1)
#44600
b10001001101010111100110111101111 E
0)
#44700
1(
1M
b100 O
0/
1)
#44800
b1 2
b1 5
0)
#44900
0K
b101 O
1)
#45000
b11 2
b11 5
0)
#45100
b10 :
b10 O
1)
#45200
0(
0M
b10010001101000101011001111 $
b10010001101000101011001111 4
b10010001101000101011001111 ;
b10011010101111001101111011110 E
0)
#45300
b1 L
b1 8
1)
#45400
b100110101011110011011110111100 E
b10 2
b10 5
b100100011010001010110011110 $
b100100011010001010110011110 4
b100100011010001010110011110 ;
0)
#45500
b10 8
b10 L
1)
#45600
b0 2
b0 5
b1001000110100010101100111100 $
b1001000110100010101100111100 4
b1001000110100010101100111100 ;
b1001101010111100110111101111000 E
0)
#45700
b11 L
b11 8
1)
#45800
1(
1M
b10011010101111001101111011110000 E
b10010001101000101011001111000 $
b10010001101000101011001111000 4
b10010001101000101011001111000 ;
0)
#45900
b100 8
b100 L
1)
#46000
0(
0M
b1 2
b1 5
b100100011010001010110011110001 $
b100100011010001010110011110001 4
b100100011010001010110011110001 ;
b110101011110011011110111100000 E
0)
#46100
b101 L
b101 8
1)
#46200
b1101010111100110111101111000000 E
b10 2
b10 5
b1001000110100010101100111100010 $
b1001000110100010101100111100010 4
b1001000110100010101100111100010 ;
0)
#46300
b110 8
b110 L
1)
#46400
1(
1M
b0 2
b0 5
b10010001101000101011001111000100 $
b10010001101000101011001111000100 4
b10010001101000101011001111000100 ;
b11010101111001101111011110000000 E
0)
#46500
b111 L
b111 8
1)
#46600
b10101011110011011110111100000000 E
b1 2
b1 5
b100011010001010110011110001001 $
b100011010001010110011110001001 4
b100011010001010110011110001001 ;
0)
#46700
b1000 8
b1000 L
1)
#46800
0(
0M
b11 2
b11 5
b1000110100010101100111100010011 $
b1000110100010101100111100010011 4
b1000110100010101100111100010011 ;
b1010111100110111101111000000000 E
0)
#46900
b1001 L
b1001 8
1)
#47000
1(
1M
b10101111001101111011110000000000 E
b10 2
b10 5
b10001101000101011001111000100110 $
b10001101000101011001111000100110 4
b10001101000101011001111000100110 ;
0)
#47100
b1010 8
b1010 L
1)
#47200
0(
0M
b1 2
b1 5
b11010001010110011110001001101 $
b11010001010110011110001001101 4
b11010001010110011110001001101 ;
b1011110011011110111100000000000 E
0)
#47300
b1011 L
b1011 8
1)
#47400
1(
1M
b10111100110111101111000000000000 E
b10 2
b10 5
b110100010101100111100010011010 $
b110100010101100111100010011010 4
b110100010101100111100010011010 ;
0)
#47500
b1100 8
b1100 L
1)
#47600
0(
0M
b1 2
b1 5
b1101000101011001111000100110101 $
b1101000101011001111000100110101 4
b1101000101011001111000100110101 ;
b1111001101111011110000000000000 E
0)
#47700
b1101 L
b1101 8
1)
#47800
1(
1M
b11110011011110111100000000000000 E
b10 2
b10 5
b11010001010110011110001001101010 $
b11010001010110011110001001101010 4
b11010001010110011110001001101010 ;
0)
#47900
b1110 8
b1110 L
1)
#48000
b1 2
b1 5
b10100010101100111100010011010101 $
b10100010101100111100010011010101 4
b10100010101100111100010011010101 ;
b11100110111101111000000000000000 E
0)
#48100
b1111 L
b1111 8
1)
#48200
b11001101111011110000000000000000 E
b11 2
b11 5
b1000101011001111000100110101011 $
b1000101011001111000100110101011 4
b1000101011001111000100110101011 ;
0)
#48300
b10000 8
b10000 L
1)
#48400
b10001010110011110001001101010111 $
b10001010110011110001001101010111 4
b10001010110011110001001101010111 ;
b10011011110111100000000000000000 E
0)
#48500
b10001 L
b10001 8
1)
#48600
0(
0M
b110111101111000000000000000000 E
b10101100111100010011010101111 $
b10101100111100010011010101111 4
b10101100111100010011010101111 ;
0)
#48700
b10010 8
b10010 L
1)
#48800
b10 2
b10 5
b101011001111000100110101011110 $
b101011001111000100110101011110 4
b101011001111000100110101011110 ;
b1101111011110000000000000000000 E
0)
#48900
b10011 L
b10011 8
1)
#49000
1(
1M
b11011110111100000000000000000000 E
b0 2
b0 5
b1010110011110001001101010111100 $
b1010110011110001001101010111100 4
b1010110011110001001101010111100 ;
0)
#49100
b10100 8
b10100 L
1)
#49200
b1 2
b1 5
b10101100111100010011010101111001 $
b10101100111100010011010101111001 4
b10101100111100010011010101111001 ;
b10111101111000000000000000000000 E
0)
#49300
b10101 L
b10101 8
1)
#49400
0(
0M
b1111011110000000000000000000000 E
b11 2
b11 5
b1011001111000100110101011110011 $
b1011001111000100110101011110011 4
b1011001111000100110101011110011 ;
0)
#49500
b10110 8
b10110 L
1)
#49600
1(
1M
b10 2
b10 5
b10110011110001001101010111100110 $
b10110011110001001101010111100110 4
b10110011110001001101010111100110 ;
b11110111100000000000000000000000 E
0)
#49700
b10111 L
b10111 8
1)
#49800
b11101111000000000000000000000000 E
b1 2
b1 5
b1100111100010011010101111001101 $
b1100111100010011010101111001101 4
b1100111100010011010101111001101 ;
0)
#49900
b11000 8
b11000 L
1)
#50000
b11 2
b11 5
b11001111000100110101011110011011 $
b11001111000100110101011110011011 4
b11001111000100110101011110011011 ;
b11011110000000000000000000000000 E
0)
#50100
b11001 L
b11001 8
1)
#50200
b10111100000000000000000000000000 E
b10011110001001101010111100110111 $
b10011110001001101010111100110111 4
b10011110001001101010111100110111 ;
0)
#50300
b11010 8
b11010 L
1)
#50400
0(
0M
b111100010011010101111001101111 $
b111100010011010101111001101111 4
b111100010011010101111001101111 ;
b1111000000000000000000000000000 E
0)
#50500
b11011 L
b11011 8
1)
#50600
1(
1M
b11110000000000000000000000000000 E
b10 2
b10 5
b1111000100110101011110011011110 $
b1111000100110101011110011011110 4
b1111000100110101011110011011110 ;
0)
#50700
b11100 8
b11100 L
1)
#50800
b1 2
b1 5
b11110001001101010111100110111101 $
b11110001001101010111100110111101 4
b11110001001101010111100110111101 ;
b11100000000000000000000000000000 E
0)
#50900
b11101 L
b11101 8
1)
#51000
b11000000000000000000000000000000 E
b11 2
b11 5
b11100010011010101111001101111011 $
b11100010011010101111001101111011 4
b11100010011010101111001101111011 ;
0)
#51100
b11110 8
b11110 L
1)
#51200
b11000100110101011110011011110111 $
b11000100110101011110011011110111 4
b11000100110101011110011011110111 ;
b10000000000000000000000000000000 E
0)
#51300
b11111 L
b11111 8
1)
#51400
0(
0M
b0 E
b10001001101010111100110111101111 $
b10001001101010111100110111101111 4
b10001001101010111100110111101111 ;
0)
#51500
b11 :
b0 8
b11 O
b0 L
1)
#51600
b10 2
b10 5
0)
#51700
1%
09
17
b1 :
1)
#51800
b0 2
b0 5
0)
#51900
1'
1>
b110 @
b0 :
1)
#52000
b1 A
b1 D
0)
#52100
0'
0>
0%
19
b111 @
1+
1)
#52200
b10 A
b10 D
0)
#52300
b0 @
07
1K
b100010010001000110011 -
b100010010001000110011 B
b100010010001000110011 Q
0+
1)
#52400
b0 A
b0 D
0)
#52500
b1 O
1)
#52600
0)
#52700
b0 O
1#
0N
1)
#52800
0)
#52900
1)
#53000
0)
#53100
0#
1N
1/
1)
#53200
b100010010001000110011 E
0)
#53300
1(
1M
b100 O
0/
1)
#53400
b1 2
b1 5
0)
#53500
b101 O
0K
1)
#53600
b11 2
b11 5
0)
#53700
0(
0M
b10 O
b10 :
1)
#53800
b1000100100010001100110 E
b10 2
b10 5
b10011010101111001101111011110 $
b10011010101111001101111011110 4
b10011010101111001101111011110 ;
0)
#53900
b1 8
b1 L
1)
#54000
b0 2
b0 5
b100110101011110011011110111100 $
b100110101011110011011110111100 4
b100110101011110011011110111100 ;
b10001001000100011001100 E
0)
#54100
b10 L
b10 8
1)
#54200
b100010010001000110011000 E
b1001101010111100110111101111000 $
b1001101010111100110111101111000 4
b1001101010111100110111101111000 ;
0)
#54300
b11 8
b11 L
1)
#54400
b10011010101111001101111011110000 $
b10011010101111001101111011110000 4
b10011010101111001101111011110000 ;
b1000100100010001100110000 E
0)
#54500
b100 L
b100 8
1)
#54600
b10001001000100011001100000 E
b110101011110011011110111100000 $
b110101011110011011110111100000 4
b110101011110011011110111100000 ;
0)
#54700
b101 8
b101 L
1)
#54800
b1101010111100110111101111000000 $
b1101010111100110111101111000000 4
b1101010111100110111101111000000 ;
b100010010001000110011000000 E
0)
#54900
b110 L
b110 8
1)
#55000
b1000100100010001100110000000 E
b11010101111001101111011110000000 $
b11010101111001101111011110000000 4
b11010101111001101111011110000000 ;
0)
#55100
b111 8
b111 L
1)
#55200
b10101011110011011110111100000000 $
b10101011110011011110111100000000 4
b10101011110011011110111100000000 ;
b10001001000100011001100000000 E
0)
#55300
b1000 L
b1000 8
1)
#55400
b100010010001000110011000000000 E
b1010111100110111101111000000000 $
b1010111100110111101111000000000 4
b1010111100110111101111000000000 ;
0)
#55500
b1001 8
b1001 L
1)
#55600
b10101111001101111011110000000000 $
b10101111001101111011110000000000 4
b10101111001101111011110000000000 ;
b1000100100010001100110000000000 E
0)
#55700
b1010 L
b1010 8
1)
#55800
1(
1M
b10001001000100011001100000000000 E
b1011110011011110111100000000000 $
b1011110011011110111100000000000 4
b1011110011011110111100000000000 ;
0)
#55900
b1011 8
b1011 L
1)
#56000
0(
0M
b1 2
b1 5
b10111100110111101111000000000001 $
b10111100110111101111000000000001 4
b10111100110111101111000000000001 ;
b10010001000110011000000000000 E
0)
#56100
b1100 L
b1100 8
1)
#56200
b100100010001100110000000000000 E
b10 2
b10 5
b1111001101111011110000000000010 $
b1111001101111011110000000000010 4
b1111001101111011110000000000010 ;
0)
#56300
b1101 8
b1101 L
1)
#56400
b0 2
b0 5
b11110011011110111100000000000100 $
b11110011011110111100000000000100 4
b11110011011110111100000000000100 ;
b1001000100011001100000000000000 E
0)
#56500
b1110 L
b1110 8
1)
#56600
1(
1M
b10010001000110011000000000000000 E
b11100110111101111000000000001000 $
b11100110111101111000000000001000 4
b11100110111101111000000000001000 ;
0)
#56700
b1111 8
b1111 L
1)
#56800
0(
0M
b1 2
b1 5
b11001101111011110000000000010001 $
b11001101111011110000000000010001 4
b11001101111011110000000000010001 ;
b100010001100110000000000000000 E
0)
#56900
b10000 L
b10000 8
1)
#57000
b1000100011001100000000000000000 E
b10 2
b10 5
b10011011110111100000000000100010 $
b10011011110111100000000000100010 4
b10011011110111100000000000100010 ;
0)
#57100
b10001 8
b10001 L
1)
#57200
1(
1M
b0 2
b0 5
b110111101111000000000001000100 $
b110111101111000000000001000100 4
b110111101111000000000001000100 ;
b10001000110011000000000000000000 E
0)
#57300
b10010 L
b10010 8
1)
#57400
0(
0M
b10001100110000000000000000000 E
b1 2
b1 5
b1101111011110000000000010001001 $
b1101111011110000000000010001001 4
b1101111011110000000000010001001 ;
0)
#57500
b10011 8
b10011 L
1)
#57600
b10 2
b10 5
b11011110111100000000000100010010 $
b11011110111100000000000100010010 4
b11011110111100000000000100010010 ;
b100011001100000000000000000000 E
0)
#57700
b10100 L
b10100 8
1)
#57800
b1000110011000000000000000000000 E
b0 2
b0 5
b10111101111000000000001000100100 $
b10111101111000000000001000100100 4
b10111101111000000000001000100100 ;
0)
#57900
b10101 8
b10101 L
1)
#58000
1(
1M
b1111011110000000000010001001000 $
b1111011110000000000010001001000 4
b1111011110000000000010001001000 ;
b10001100110000000000000000000000 E
0)
#58100
b10110 L
b10110 8
1)
#58200
0(
0M
b11001100000000000000000000000 E
b1 2
b1 5
b11110111100000000000100010010001 $
b11110111100000000000100010010001 4
b11110111100000000000100010010001 ;
0)
#58300
b10111 8
b10111 L
1)
#58400
b10 2
b10 5
b11101111000000000001000100100010 $
b11101111000000000001000100100010 4
b11101111000000000001000100100010 ;
b110011000000000000000000000000 E
0)
#58500
b11000 L
b11000 8
1)
#58600
b1100110000000000000000000000000 E
b0 2
b0 5
b11011110000000000010001001000100 $
b11011110000000000010001001000100 4
b11011110000000000010001001000100 ;
0)
#58700
b11001 8
b11001 L
1)
#58800
1(
1M
b10111100000000000100010010001000 $
b10111100000000000100010010001000 4
b10111100000000000100010010001000 ;
b11001100000000000000000000000000 E
0)
#58900
b11010 L
b11010 8
1)
#59000
b10011000000000000000000000000000 E
b1 2
b1 5
b1111000000000001000100100010001 $
b1111000000000001000100100010001 4
b1111000000000001000100100010001 ;
0)
#59100
b11011 8
b11011 L
1)
#59200
0(
0M
b11 2
b11 5
b11110000000000010001001000100011 $
b11110000000000010001001000100011 4
b11110000000000010001001000100011 ;
b110000000000000000000000000000 E
0)
#59300
b11100 L
b11100 8
1)
#59400
b1100000000000000000000000000000 E
b10 2
b10 5
b11100000000000100010010001000110 $
b11100000000000100010010001000110 4
b11100000000000100010010001000110 ;
0)
#59500
b11101 8
b11101 L
1)
#59600
1(
1M
b0 2
b0 5
b11000000000001000100100010001100 $
b11000000000001000100100010001100 4
b11000000000001000100100010001100 ;
b11000000000000000000000000000000 E
0)
#59700
b11110 L
b11110 8
1)
#59800
b10000000000000000000000000000000 E
b1 2
b1 5
b10000000000010001001000100011001 $
b10000000000010001001000100011001 4
b10000000000010001001000100011001 ;
0)
#59900
b11111 8
b11111 L
1)
#60000
0(
0M
b11 2
b11 5
b100010010001000110011 $
b100010010001000110011 4
b100010010001000110011 ;
b0 E
0)
#60100
b0 L
b11 O
b0 8
b11 :
1)
#60200
b10 2
b10 5
0)
#60300
b1 :
17
1%
09
1)
#60400
b0 2
b0 5
0)
#60500
1'
1>
b0 :
b110 @
1)
#60600
b1 A
b1 D
0)
#60700
0'
0>
b111 @
0%
19
1+
1)
#60800
b10 A
b10 D
0)
#60900
1K
07
b0 @
b1000100010101010110011001110111 -
b1000100010101010110011001110111 B
b1000100010101010110011001110111 Q
0+
1)
#61000
b0 A
b0 D
0)
#61100
b1 O
1)
#61200
0)
#61300
1#
0N
b0 O
1)
#61400
0)
#61500
1)
#61600
0)
#61700
0#
1N
1/
1)
#61800
b1000100010101010110011001110111 E
0)
#61900
1(
1M
b100 O
0/
1)
#62000
b1 2
b1 5
0)
#62100
0K
b101 O
1)
#62200
b11 2
b11 5
0)
#62300
0(
0M
b10 :
b10 O
1)
#62400
1(
1M
b10 2
b10 5
b1000100100010001100110 $
b1000100100010001100110 4
b1000100100010001100110 ;
b10001000101010101100110011101110 E
0)
#62500
b1 L
b1 8
1)
#62600
0(
0M
b10001010101011001100111011100 E
b1 2
b1 5
b10001001000100011001101 $
b10001001000100011001101 4
b10001001000100011001101 ;
0)
#62700
b10 8
b10 L
1)
#62800
b10 2
b10 5
b100010010001000110011010 $
b100010010001000110011010 4
b100010010001000110011010 ;
b100010101010110011001110111000 E
0)
#62900
b11 L
b11 8
1)
#63000
b1000101010101100110011101110000 E
b0 2
b0 5
b1000100100010001100110100 $
b1000100100010001100110100 4
b1000100100010001100110100 ;
0)
#63100
b100 8
b100 L
1)
#63200
1(
1M
b10001001000100011001101000 $
b10001001000100011001101000 4
b10001001000100011001101000 ;
b10001010101011001100111011100000 E
0)
#63300
b101 L
b101 8
1)
#63400
0(
0M
b10101010110011001110111000000 E
b1 2
b1 5
b100010010001000110011010001 $
b100010010001000110011010001 4
b100010010001000110011010001 ;
0)
#63500
b110 8
b110 L
1)
#63600
b10 2
b10 5
b1000100100010001100110100010 $
b1000100100010001100110100010 4
b1000100100010001100110100010 ;
b101010101100110011101110000000 E
0)
#63700
b111 L
b111 8
1)
#63800
b1010101011001100111011100000000 E
b0 2
b0 5
b10001001000100011001101000100 $
b10001001000100011001101000100 4
b10001001000100011001101000100 ;
0)
#63900
b1000 8
b1000 L
1)
#64000
1(
1M
b100010010001000110011010001000 $
b100010010001000110011010001000 4
b100010010001000110011010001000 ;
b10101010110011001110111000000000 E
0)
#64100
b1001 L
b1001 8
1)
#64200
0(
0M
b1010101100110011101110000000000 E
b1 2
b1 5
b1000100100010001100110100010001 $
b1000100100010001100110100010001 4
b1000100100010001100110100010001 ;
0)
#64300
b1010 8
b1010 L
1)
#64400
1(
1M
b10 2
b10 5
b10001001000100011001101000100010 $
b10001001000100011001101000100010 4
b10001001000100011001101000100010 ;
b10101011001100111011100000000000 E
0)
#64500
b1011 L
b1011 8
1)
#64600
0(
0M
b1010110011001110111000000000000 E
b1 2
b1 5
b10010001000110011010001000101 $
b10010001000110011010001000101 4
b10010001000110011010001000101 ;
0)
#64700
b1100 8
b1100 L
1)
#64800
1(
1M
b10 2
b10 5
b100100010001100110100010001010 $
b100100010001100110100010001010 4
b100100010001100110100010001010 ;
b10101100110011101110000000000000 E
0)
#64900
b1101 L
b1101 8
1)
#65000
0(
0M
b1011001100111011100000000000000 E
b1 2
b1 5
b1001000100011001101000100010101 $
b1001000100011001101000100010101 4
b1001000100011001101000100010101 ;
0)
#65100
b1110 8
b1110 L
1)
#65200
1(
1M
b10 2
b10 5
b10010001000110011010001000101010 $
b10010001000110011010001000101010 4
b10010001000110011010001000101010 ;
b10110011001110111000000000000000 E
0)
#65300
b1111 L
b1111 8
1)
#65400
0(
0M
b1100110011101110000000000000000 E
b1 2
b1 5
b100010001100110100010001010101 $
b100010001100110100010001010101 4
b100010001100110100010001010101 ;
0)
#65500
b10000 8
b10000 L
1)
#65600
1(
1M
b10 2
b10 5
b1000100011001101000100010101010 $
b1000100011001101000100010101010 4
b1000100011001101000100010101010 ;
b11001100111011100000000000000000 E
0)
#65700
b10001 L
b10001 8
1)
#65800
b10011001110111000000000000000000 E
b1 2
b1 5
b10001000110011010001000101010101 $
b10001000110011010001000101010101 4
b10001000110011010001000101010101 ;
0)
#65900
b10010 8
b10010 L
1)
#66000
0(
0M
b11 2
b11 5
b10001100110100010001010101011 $
b10001100110100010001010101011 4
b10001100110100010001010101011 ;
b110011101110000000000000000000 E
0)
#66100
b10011 L
b10011 8
1)
#66200
b1100111011100000000000000000000 E
b10 2
b10 5
b100011001101000100010101010110 $
b100011001101000100010101010110 4
b100011001101000100010101010110 ;
0)
#66300
b10100 8
b10100 L
1)
#66400
1(
1M
b0 2
b0 5
b1000110011010001000101010101100 $
b1000110011010001000101010101100 4
b1000110011010001000101010101100 ;
b11001110111000000000000000000000 E
0)
#66500
b10101 L
b10101 8
1)
#66600
b10011101110000000000000000000000 E
b1 2
b1 5
b10001100110100010001010101011001 $
b10001100110100010001010101011001 4
b10001100110100010001010101011001 ;
0)
#66700
b10110 8
b10110 L
1)
#66800
0(
0M
b11 2
b11 5
b11001101000100010101010110011 $
b11001101000100010101010110011 4
b11001101000100010101010110011 ;
b111011100000000000000000000000 E
0)
#66900
b10111 L
b10111 8
1)
#67000
b1110111000000000000000000000000 E
b10 2
b10 5
b110011010001000101010101100110 $
b110011010001000101010101100110 4
b110011010001000101010101100110 ;
0)
#67100
b11000 8
b11000 L
1)
#67200
1(
1M
b0 2
b0 5
b1100110100010001010101011001100 $
b1100110100010001010101011001100 4
b1100110100010001010101011001100 ;
b11101110000000000000000000000000 E
0)
#67300
b11001 L
b11001 8
1)
#67400
b11011100000000000000000000000000 E
b1 2
b1 5
b11001101000100010101010110011001 $
b11001101000100010101010110011001 4
b11001101000100010101010110011001 ;
0)
#67500
b11010 8
b11010 L
1)
#67600
b11 2
b11 5
b10011010001000101010101100110011 $
b10011010001000101010101100110011 4
b10011010001000101010101100110011 ;
b10111000000000000000000000000000 E
0)
#67700
b11011 L
b11011 8
1)
#67800
0(
0M
b1110000000000000000000000000000 E
b110100010001010101011001100111 $
b110100010001010101011001100111 4
b110100010001010101011001100111 ;
0)
#67900
b11100 8
b11100 L
1)
#68000
1(
1M
b10 2
b10 5
b1101000100010101010110011001110 $
b1101000100010101010110011001110 4
b1101000100010101010110011001110 ;
b11100000000000000000000000000000 E
0)
#68100
b11101 L
b11101 8
1)
#68200
b11000000000000000000000000000000 E
b1 2
b1 5
b11010001000101010101100110011101 $
b11010001000101010101100110011101 4
b11010001000101010101100110011101 ;
0)
#68300
b11110 8
b11110 L
1)
#68400
b11 2
b11 5
b10100010001010101011001100111011 $
b10100010001010101011001100111011 4
b10100010001010101011001100111011 ;
b10000000000000000000000000000000 E
0)
#68500
b11111 L
b11111 8
1)
#68600
0(
0M
b0 E
b1000100010101010110011001110111 $
b1000100010101010110011001110111 4
b1000100010101010110011001110111 ;
0)
#68700
b11 :
b0 8
b11 O
b0 L
1)
#68800
b10 2
b10 5
0)
#68900
1%
09
17
b1 :
1)
#69000
b0 2
b0 5
0)
#69100
1'
1>
b110 @
b0 :
1)
#69200
b1 A
b1 D
0)
#69300
0'
0>
0%
19
b111 @
1+
1)
#69400
b10 A
b10 D
0)
#69500
b0 @
07
1K
0+
1)
#69600
b0 A
b0 D
0)
#69700
b1 O
1)
#69800
0)
#69900
b0 O
1#
0N
1)
#70000
0)
#70100
1)
#70200
0)
#70300
1)
#70400
0)
#70500
1)
#70600
0)
#70700
1)
#70800
0)
#70900
1)
#71000
0)
#71100
1)
#71200
0)
#71300
1)
#71400
0)
#71500
1)
#71600
0)
#71700
1)
#71800
0)
#71900
1)
#72000
0)
#72100
1)
#72200
0)
#72300
1)
#72400
0)
#72500
1)
#72600
0)
#72700
1)
#72800
0)
#72900
1)
#73000
0)
#73100
1)
#73200
0)
#73300
1)
#73400
0)
#73500
1)
#73600
0)
#73700
1)
#73800
0)
#73900
1)
#74000
0)
#74100
1)
#74200
0)
#74300
1)
#74400
0)
#74500
1)
#74600
0)
#74700
1)
#74800
0)
#74900
1)
#75000
0)
#75100
1)
#75200
0)
#75300
1)
#75400
0)
#75500
1)
#75600
0)
#75700
1)
#75800
0)
#75900
1)
#76000
0)
#76100
1)
#76200
0)
#76300
1)
#76400
0)
#76500
1)
#76600
0)
#76700
1)
#76800
0)
#76900
1)
#77000
0)
#77100
1)
#77200
0)
#77300
1)
#77400
0)
#77500
1)
#77600
0)
#77700
1)
#77800
0)
#77900
1)
#78000
0)
#78100
1)
#78200
0)
#78300
1)
#78400
0)
#78500
1)
#78600
0)
#78700
1)
#78800
0)
#78900
1)
#79000
0)
#79100
1)
#79200
0)
#79300
1)
#79400
0)
#79500
1)
